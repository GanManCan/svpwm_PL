----------------------------------------------------------------------------
--  % Name        : svpwm_pl_tb_pkg.vhdl %                                   --
--  % Project     :    %                                   --
--  % Version     : 1.0               %                                   --
--  % Created_By  :     %                                   --
--  % Date_Created: 2022-02-12        %                                   --
--                                                                        --
--  Description:                                                          --
--                                                                        --
----------------------------------------------------------------------------
--  Revision History                                                      --
--                                                                        --
--  Version    Date       Sign       Change Description                   --
--  ------- ----------  ----------   ------------------                   --
--                       --
--                                                                        --
----------------------------------------------------------------------------
--  TODO List                                                             --
--                                                                        -- 
--                                                                        --
----------------------------------------------------------------------------

----------------------------------------------------------------------------
-- Configuration Declaration.
----------------------------------------------------------------------------

----------------------------------------------------------------------------
-- Library Declaration.
----------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


----------------------------------------------------------------------------
-- PACKAGE DECLARATION.
----------------------------------------------------------------------------
PACKAGE svpwm_pl_tb_pkg IS
----------------------------------------------------------------------------
-- Global Constant Declaration.  
----------------------------------------------------------------------------


----------------------------------------------------------------------------
-- Procedures Declaration.  
----------------------------------------------------------------------------
  PROCEDURE pulse_high(SIGNAL clk    : IN  STD_LOGIC;
                       SIGNAL pulsed : OUT STD_LOGIC);

                          

END PACKAGE svpwm_pl_tb_pkg;


----------------------------------------------------------------------------
-- PACKAGE BODY DECLARATION.
----------------------------------------------------------------------------
PACKAGE BODY svpwm_pl_tb_pkg is

----------------------------------------------------------------------------
-- Procedures Implementation.  
----------------------------------------------------------------------------
  PROCEDURE pulse_high(SIGNAL clk    : IN  STD_LOGIC;
                       SIGNAL pulsed : OUT STD_LOGIC) IS
  BEGIN
    pulsed <= '1';
    WAIT UNTIL rising_edge(clk);
    pulsed <= '0';
  END PROCEDURE pulse_high;

  
END PACKAGE BODY svpwm_pl_tb_pkg;
